module pc (
	input logic 		clk,
	input logic 		rst,
	input logic [31:0] 	pc_i,
	output logic [31:0] pc_o
);

endmodule
