module mux_a (
    input logic [31:0] pc_o,
    input logic [31:0] rs1_data
);

endmodule