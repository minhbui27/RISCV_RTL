module main_ctrl (
    input  logic [31:0] inst,
    output logic        reg_wr,
    output logic [3:0]  alu_op,
    output logic        sel_a,
    output logic        sel_b,
    output logic        mem_wr,
    output logic        mem_rd,
    output logic [2:0]  mask,
    output logic [1:0]  sel_wb

);

endmodule