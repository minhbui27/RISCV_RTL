`timescale 1ns/1ns
module mux_wb (
    input logic [31:0] dmem_o,
    input logic [31:0] pc_p4,
    input logic [31:0] alu_o
);


endmodule
