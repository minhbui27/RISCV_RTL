module mux_b (
    input logic [31:0] rs2_data,
    input logic [31:0] imm_o
);

endmodule