`timescale 1ns/1ns
module imm_gen (
	input [31:0]	inst,
	output [31:0] 	imm_o
);

endmodule
